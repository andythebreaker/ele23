** Profile: "Example PS.6.2 Rout-AC"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.6\appendix b-ps.6-example ps.6.2 rout-ac.sim ] 

** Creating circuit file "appendix b-ps.6-example ps.6.2 rout-ac.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 25 0.1 100E6
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.6.2 Rout.net"


.END
