** Profile: "Example PS.2.2 AC Gain-AC2"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\CHAPTER 2\Appendix B-PS.2-Example PS.2.2 AC Gain-AC2.sim ] 

** Creating circuit file "Appendix B-PS.2-Example PS.2.2 AC Gain-AC2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "..\sedra_lib.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 25 1 10E6
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\Appendix B-PS.2-Example PS.2.2 AC Gain.net" 


.END
