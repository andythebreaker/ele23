** Profile: "Example PS.9.1-Bias"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.9\appendix b-ps.9-example ps.9.1-bias.sim ] 

** Creating circuit file "appendix b-ps.9-example ps.9.1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "../Example PS.9.1.net"


.END
