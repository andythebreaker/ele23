** Profile: "Example PS.2.1 Step Response-Transient"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\CHAPTER 2\appendix b-ps.2-example ps.2.1 step response-transient.sim ] 

** Creating circuit file "appendix b-ps.2-example ps.2.1 step response-transient.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 140us 0 10n 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.2.1 Step Response.net"


.END
