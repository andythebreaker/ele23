** Profile: "Example PS.2.2 Slew Rate-Transient"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\CHAPTER 2\appendix b-ps.2-example ps.2.2 slew rate-transient.sim ] 

** Creating circuit file "appendix b-ps.2-example ps.2.2 slew rate-transient.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80u 0 10n 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.2.2 Slew Rate.net"


.END
