** Profile: "Example 9.4 Opamp-DC Transfer"  [ C:\Documents and Settings\Adel Sedra\My Documents\SEDRA WORK\SEDRA-PSPICE-CD\CHAPTER 9\chapter 9-Example 9.4 Opamp-DC Transfer.sim ] 

** Creating circuit file "chapter 9-Example 9.4 Opamp-DC Transfer.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "..\sedra_lib.lib" 
* From [PSPICE NETLIST] section of e:\cadence\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_Vd -5m 5m 1u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\chapter 9-Example 9.4 Opamp.net" 


.END
