** Profile: "Example PS.5.1 AC Gain-AC"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.5\appendix b-ps.5-example ps.5.1 ac gain-ac.sim ] 

** Creating circuit file "appendix b-ps.5-example ps.5.1 ac gain-ac.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 25 0.0001 1E10
.STEP PARAM CS LIST 1E-15 10u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.5.1 AC Gain.net"


.END
