** Profile: "zener test-DC Sweep"  [ C:\Documents and Settings\Adel Sedra\My Documents\SEDRA WORK\PSPICE Archive\CHAPTER 3\chapter 3-zener test-DC Sweep.sim ] 

** Creating circuit file "chapter 3-zener test-DC Sweep.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:\Documents and Settings\Adel Sedra\My Documents\SEDRA WORK\PSPICE Libraries\sedra_lib.lib" 
* From [PSPICE NETLIST] section of e:\cadence\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_Vtest 0 6 1m 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\chapter 3-zener test.net" 


.END
