** Profile: "Example PS.12.1 Slew Rate-slew"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.12\appendix b-ps.12-example ps.12.1 slew rate-slew.sim ] 

** Creating circuit file "appendix b-ps.12-example ps.12.1 slew rate-slew.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.25u 0 0.01n 
.STEP PARAM R LIST 1.53K 3.2K 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.12.1 Slew Rate.net"


.END
