** Profile: "Example PS.12.1 AC Gain-AC"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.12\appendix b-ps.12-example ps.12.1 ac gain-ac.sim ] 

** Creating circuit file "appendix b-ps.12-example ps.12.1 ac gain-ac.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 20 1 10E9
.STEP PARAM Cc LIST 1E-15 0.6p 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.12.1 AC Gain.net"


.END
