** Profile: "Example PS.4.1-transient"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.4\appendix b-ps.4-example ps.4.1-transient.sim ] 

** Creating circuit file "appendix b-ps.4-example ps.4.1-transient.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 200m 0 20u 
.STEP PARAM Rload LIST 150 200 250 500 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC "../Example PS.4.1.net"


.END
