** Profile: "Class B Output Stage-Transient"  [ C:\Documents and Settings\Adel Sedra\My Documents\SEDRA WORK\SEDRA-PSPICE-CD\CHAPTER 14\chapter 14-Class B Output Stage-Transient.sim ] 

** Creating circuit file "chapter 14-Class B Output Stage-Transient.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "..\sedra_lib.lib" 
* From [PSPICE NETLIST] section of e:\cadence\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 10u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\chapter 14-Class B Output Stage.net" 


.END
