** Profile: "CMOS Opamp-AC"  [ C:\Documents and Settings\Adel Sedra\My Documents\SEDRA WORK\SEDRA-PSPICE-CD\CHAPTER 9\chapter 9-CMOS Opamp-AC.sim ] 

** Creating circuit file "chapter 9-CMOS Opamp-AC.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "..\sedra_lib.lib" 
* From [PSPICE NETLIST] section of e:\cadence\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 20 1 10E9
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\chapter 9-CMOS Opamp.net" 


.END
