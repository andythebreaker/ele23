** Profile: "Example PS.9.1-DC Sweep"  [ C:\Users\Behrooz\Desktop\SPICE Examples\Appendix B-PS.9\appendix b-ps.9-example ps.9.1-dc sweep.sim ] 

** Creating circuit file "Appendix B-PS.9-Example PS.9.1-DC Sweep.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\OrCAD\OrCAD_16.0\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_Vin 1 2.5 0.1m 
.STEP PARAM W LIST 10.65u 12.5u 14.37u 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.9.1.net"


.END
