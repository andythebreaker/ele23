** Profile: "Example PS.8.1-Differential DC Transfer"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\Appendix B-PS.8\appendix b-ps.8-example ps.8.1-differential dc transfer.sim ] 

** Creating circuit file "appendix b-ps.8-example ps.8.1-differential dc transfer.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "C:/Users/Behrooz/Desktop/SPICE Examples - Orcad New Version/sedra_lib.lib"
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_Vd -5m 5m 0.001m 
.STEP PARAM R3_2 LIST 0.00001 3K 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "../Example PS.8.1.net"


.END
