** Profile: "Example PS.2.1 Rout-Example PS.2.1 Rout-AC1"  [ C:\Documents and Settings\Administrator\My Documents\SPICE Examples Converted\CHAPTER 2\appendix b-ps.2-example ps.2.1 rout-example ps.2.1 rout-ac1.sim ] 

** Creating circuit file "appendix b-ps.2-example ps.2.1 rout-example ps.2.1 rout-ac1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.LIB "..\sedra_lib.lib" 
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 25 0.1 100E6
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC ".\Appendix B-PS.2-Example PS.2.1 Rout.net" 


.END
